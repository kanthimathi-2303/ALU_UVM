//`ifndef DEFINES_V
//`define DEFINES_V

`define DATA_WIDTH 8
`define CMD_WIDTH 4
`define NO_OF_TRANS 10

//`endif
